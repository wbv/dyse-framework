--| test_pad: a scratchpad for testing small pieces of VHDL
--|

library ieee;
use ieee.std_logic_1164.all;

entity test_pad is
end test_pad;

architecture behavioral of test_pad is
begin
end behavioral;
