../vivado/ip/count_stream_test_0.1/hdl/count_stream_test_v0_1_S_AXI_registers.vhd